-------------------------------------------------------------------------
-- Will Galles
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------


-- tb_reg_N.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains a simple VHDL testbench for the
-- edge-triggered flip-flop with parallel access and reset.
--
--
-- NOTES:
-- 8/19/16 by JAZ::Design created.
-- 11/25/19 by H3:Changed name to avoid name conflict with Quartus
--          primitives.
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_reg_N is
  generic(gCLK_HPER   : time := 50 ns);
end tb_reg_N;

architecture behavior of tb_reg_N is
  
  -- Calculate the clock period as twice the half-period
  constant cCLK_PER  : time := gCLK_HPER * 2;
  constant n : integer :=16;

  component reg_N
    generic(N : integer := 16);
    port(i_CLK        : in std_logic;     -- Clock input
         i_RST        : in std_logic;     -- Reset input
         i_WE         : in std_logic;     -- Write enable input
         i_D          : in std_logic_vector(N-1 downto 0);     -- Data value input
         o_Q          : out std_logic_vector(N-1 downto 0));   -- Data value output
  end component;

  -- Temporary signals to connect to the dff component.
  signal s_CLK, s_RST, s_WE  : std_logic;
  signal s_Q : std_logic_vector(n-1 downto 0);-- := x"0001";
  signal s_D : std_logic_vector(n-1 downto 0) := x"0000";

begin

  DUT: reg_N 
  generic map(n)
  port map(i_CLK => s_CLK, 
           i_RST => s_RST,
           i_WE  => s_WE,
           i_D   => s_D,
           o_Q   => s_Q);

  -- This process sets the clock value (low for gCLK_HPER, then high
  -- for gCLK_HPER). Absent a "wait" command, processes restart 
  -- at the beginning once they have reached the final statement.
  P_CLK: process
  begin
    s_CLK <= '0';
    wait for gCLK_HPER;
    s_CLK <= '1';
    wait for gCLK_HPER;
  end process;
  
  -- Testbench process  
  P_TB: process
  begin
    -- Reset the FF
    s_RST <= '1';
    s_WE  <= '0';
    s_D   <= x"0000";
    wait for cCLK_PER;

    -- Store '1'
    s_RST <= '0';
    s_WE  <= '1';
    s_D   <= x"0001";
    wait for cCLK_PER;  

    -- Keep '1'
    s_RST <= '0';
    s_WE  <= '0';
    s_D   <= x"0000";
    wait for cCLK_PER;  

    -- Store '0xFFFF'    
    s_RST <= '0';
    s_WE  <= '1';
    s_D   <= x"FFFF";
    wait for cCLK_PER;  

    -- Keep '0xFFFF'
    s_RST <= '0';
    s_WE  <= '0';
    s_D   <= x"0001";
    wait for cCLK_PER;  

    -- Store '0xF007'    
    s_RST <= '0';
    s_WE  <= '1';
    s_D   <= x"F007";
    wait for cCLK_PER;  

    -- Keep 'DEAD'
    s_RST <= '0';
    s_WE  <= '0';
    s_D   <= x"DEAD";
    wait for cCLK_PER;  

    wait;
  end process;
  
end behavior;
