    Mac OS X            	   2  J     |                                      ATTR      |   �   �                  �     com.apple.lastuseddate#PS       �   H  com.apple.macl     4   H  com.apple.quarantine �u�a    ��3     �; $�J���3Rh��                                                      q/0081;61e5cbce;Microsoft\x20Teams;B65EF45D-A64C-430E-A13E-AF746065E802 