    Mac OS X            	   2   �      �                                      ATTR       �   �   H                  �   H  com.apple.quarantine q/0081;61e5cbce;Microsoft\x20Teams;B65EF45D-A64C-430E-A13E-AF746065E802 